module c880(N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68,
     N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96,
     N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146,
     N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195,
     N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261,
     N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422,
     N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864,
     N865, N866, N874, N878, N879, N880);
  input N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72,
       N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96,
       N101, N106, N111, N116, N121, N126, N130, N135, N138, N143,
       N146, N149, N152, N153, N156, N159, N165, N171, N177, N183,
       N189, N195, N201, N207, N210, N219, N228, N237, N246, N255,
       N259, N260, N261, N267, N268;
  output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423,
       N446, N447, N448, N449, N450, N767, N768, N850, N863, N864,
       N865, N866, N874, N878, N879, N880;
  wire N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72,
       N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96,
       N101, N106, N111, N116, N121, N126, N130, N135, N138, N143,
       N146, N149, N152, N153, N156, N159, N165, N171, N177, N183,
       N189, N195, N201, N207, N210, N219, N228, N237, N246, N255,
       N259, N260, N261, N267, N268;
  wire N388, N389, N390, N391, N418, N419, N420, N421, N422, N423,
       N446, N447, N448, N449, N450, N767, N768, N850, N863, N864,
       N865, N866, N874, N878, N879, N880;
  wire N269, N270, N279, N280, N285, N287, N293, N294;
  wire N295, N296, N298, N301, N302, N303, N304, N305;
  wire N306, N307, N308, N309, N316, N317, N318, N319;
  wire N322, N323, N324, N325, N326, N327, N328, N329;
  wire N330, N331, N332, N333, N334, N335, N336, N337;
  wire N338, N339, N340, N341, N343, N347, N349, N350;
  wire N352, N355, N357, N360, N363, N366, N375, N376;
  wire N379, N382, N385, N400, N404, N405, N406, N407;
  wire N408, N409, N410, N411, N412, N413, N414, N415;
  wire N416, N417, N425, N426, N427, N442, N443, N444;
  wire N445, N460, N463, N466, N475, N476, N477, N479;
  wire N481, N483, N488, N492, N495, N498, N499, N500;
  wire N501, N502, N503, N504, N505, N506, N507, N508;
  wire N509, N510, N511, N512, N513, N514, N515, N516;
  wire N517, N518, N519, N520, N521, N522, N523, N524;
  wire N525, N526, N527, N528, N529, N530, N533, N536;
  wire N537, N538, N539, N540, N541, N542, N543, N544;
  wire N547, N550, N551, N552, N553, N557, N561, N565;
  wire N569, N573, N577, N581, N585, N586, N587, N588;
  wire N589, N590, N593, N596, N597, N600, N605, N606;
  wire N609, N615, N616, N619, N624, N625, N628, N631;
  wire N632, N635, N640, N641, N644, N650, N651, N654;
  wire N659, N662, N665, N669, N670, N673, N677, N678;
  wire N682, N686, N687, N692, N696, N697, N700, N704;
  wire N705, N708, N712, N713, N717, N721, N722, N727;
  wire N731, N732, N733, N734, N736, N737, N739, N740;
  wire N742, N743, N745, N746, N748, N749, N751, N752;
  wire N754, N755, N757, N758, N759, N760, N761, N762;
  wire N763, N764, N765, N766, N769, N770, N771, N772;
  wire N773, N777, N778, N781, N782, N785, N786, N787;
  wire N788, N789, N790, N791, N792, N793, N794, N795;
  wire N796, N802, N803, N804, N805, N806, N807, N808;
  wire N809, N810, N812, N813, N814, N815, N819, N822;
  wire N825, N826, N827, N828, N830, N831, N832, N833;
  wire N834, N835, N836, N841, N842, N843, N844, N845;
  wire N849, N851, N852, N853, N859, N860, N861, n_87;
  wire n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95;
  wire n_96;
  and AND2_18 (N391, N85, N86);
  and AND2_28 (N309, N8, N138);
  and AND2_30 (N316, N51, N138);
  and AND2_31 (N317, N17, N138);
  and AND2_32 (N318, N152, N138);
  and AND2_35 (N323, N17, N42);
  and AND2_44 (N332, N210, N91);
  and AND2_45 (N333, N210, N96);
  and AND2_46 (N334, N210, N101);
  and AND2_47 (N335, N210, N106);
  and AND2_48 (N336, N210, N111);
  and AND2_49 (N337, N255, N259);
  and AND2_50 (N338, N210, N116);
  and AND2_51 (N339, N255, N260);
  and AND2_52 (N340, N210, N121);
  and AND2_53 (N341, N255, N267);
  and AND2_68 (N423, N90, N298);
  and AND2_92 (N406, N357, N360);
  and AND2_95 (N409, N363, N366);
  and AND2_99 (N413, N376, N379);
  and AND2_102 (N416, N382, N385);
  and AND2_103 (N417, N210, N268);
  and AND2_111 (N425, N404, N405);
  and AND2_112 (N426, N407, N408);
  and AND2_118 (N444, N411, N412);
  and AND2_119 (N445, N414, N415);
  and AND2_129 (N475, N143, N427);
  and AND2_131 (N477, N146, N427);
  and AND2_133 (N479, N149, N427);
  and AND2_135 (N481, N153, N427);
  and AND2_148 (N502, N91, N466);
  and AND2_150 (N504, N96, N466);
  and AND2_152 (N506, N101, N466);
  and AND2_154 (N508, N106, N466);
  and AND2_156 (N510, N143, N483);
  and AND2_157 (N511, N111, N466);
  and AND2_158 (N512, N146, N483);
  and AND2_159 (N513, N116, N466);
  and AND2_160 (N514, N149, N483);
  and AND2_161 (N515, N121, N466);
  and AND2_162 (N516, N153, N483);
  and AND2_163 (N517, N126, N466);
  and AND2_168 (N522, N400, N159);
  and AND2_169 (N523, N400, N165);
  and AND2_170 (N524, N400, N171);
  and AND2_171 (N525, N400, N177);
  and AND2_172 (N526, N400, N183);
  and AND2_190 (N552, N530, N533);
  and AND2_201 (N587, N544, N547);
  and AND2_202 (N588, N550, N551);
  and AND2_203 (N589, N585, N586);
  and AND2_206 (N596, N246, N553);
  and AND2_209 (N605, N246, N557);
  and AND2_212 (N615, N246, N561);
  and AND2_215 (N624, N246, N565);
  and AND2_218 (N631, N246, N569);
  and AND2_221 (N640, N246, N573);
  and AND2_224 (N650, N246, N577);
  and AND2_227 (N659, N246, N581);
  and AND2_231 (N665, N593, N590);
  and AND2_234 (N673, N600, N597);
  and AND2_237 (N682, N609, N606);
  and AND2_240 (N692, N619, N616);
  and AND2_243 (N700, N628, N625);
  and AND2_246 (N708, N635, N632);
  and AND2_249 (N717, N644, N641);
  and AND2_252 (N727, N654, N651);
  and AND2_258 (N736, N228, N665);
  and AND2_259 (N737, N237, N662);
  and AND2_261 (N739, N228, N673);
  and AND2_262 (N740, N237, N670);
  and AND2_264 (N742, N228, N682);
  and AND2_265 (N743, N237, N678);
  and AND2_267 (N745, N228, N692);
  and AND2_268 (N746, N237, N687);
  and AND2_270 (N748, N228, N700);
  and AND2_271 (N749, N237, N697);
  and AND2_273 (N751, N228, N708);
  and AND2_274 (N752, N237, N705);
  and AND2_276 (N754, N228, N717);
  and AND2_277 (N755, N237, N713);
  and AND2_280 (N758, N727, N261);
  and AND2_281 (N759, N228, N727);
  and AND2_282 (N760, N237, N722);
  and AND2_304 (N789, N700, N773);
  and AND2_306 (N791, N708, N778);
  and AND2_308 (N793, N717, N782);
  and AND2_309 (N794, N219, N786);
  and AND2_317 (N807, N692, N796);
  and AND2_318 (N808, N219, N802);
  and AND2_319 (N809, N219, N803);
  and AND2_320 (N810, N219, N804);
  and AND2_334 (N831, N665, N815);
  and AND2_336 (N833, N673, N819);
  and AND2_338 (N835, N682, N822);
  and AND2_339 (N836, N219, N825);
  and AND2_352 (N849, N590, N841);
  and AND2_354 (N851, N219, N842);
  and AND2_355 (N852, N219, N843);
  and AND2_356 (N853, N219, N844);
  and AND3_3 (N390, N29, N36, N42);
  and AND3_4 (N447, N1, N26, N51);
  and AND3_10 (N287, N29, N75, N80);
  and AND3_11 (N388, N29, N75, N42);
  and AND3_12 (N389, N29, N36, N80);
  and AND3_14 (N293, N59, N75, N80);
  and AND3_15 (N294, N59, N75, N42);
  and AND3_16 (N295, N59, N36, N80);
  and AND3_17 (N296, N59, N36, N42);
  and AND3_113 (N427, N319, N447, N55);
  nand NAND2_8 (N285, N29, N68);
  nand NAND2_20 (N301, N91, N96);
  nand NAND2_22 (N303, N101, N106);
  nand NAND2_24 (N305, N111, N116);
  nand NAND2_26 (N307, N121, N126);
  nand NAND2_33 (N319, N59, N156);
  nand NAND2_36 (N324, N159, N165);
  nand NAND2_38 (N326, N171, N177);
  nand NAND2_40 (N328, N183, N189);
  nand NAND2_42 (N330, N195, N201);
  nand NAND2_67 (N355, N89, N298);
  nand NAND2_69 (N357, N301, N302);
  nand NAND2_70 (N360, N303, N304);
  nand NAND2_71 (N363, N305, N306);
  nand NAND2_72 (N366, N307, N308);
  nand NAND2_75 (N376, N324, N325);
  nand NAND2_76 (N379, N326, N327);
  nand NAND2_77 (N382, N328, N329);
  nand NAND2_78 (N385, N330, N331);
  nand NAND2_96 (N410, N347, N352);
  nand NAND2_128 (N466, N442, N410);
  nand NAND2_137 (N483, N443, N1);
  nand NAND2_144 (N498, N130, N460);
  nand NAND2_146 (N500, N463, N135);
  nand NAND2_164 (N518, N130, N492);
  nand NAND2_166 (N520, N495, N207);
  nand NAND2_173 (N527, N400, N189);
  nand NAND2_174 (N528, N400, N195);
  nand NAND2_175 (N529, N400, N201);
  nand NAND2_176 (N530, N498, N499);
  nand NAND2_177 (N533, N500, N501);
  nand NAND2_186 (N544, N518, N519);
  nand NAND2_187 (N547, N520, N521);
  nand NAND2_191 (N553, N536, N503);
  nand NAND2_192 (N557, N537, N505);
  nand NAND2_193 (N561, N538, N507);
  nand NAND2_194 (N565, N539, N509);
  nand NAND2_195 (N569, N488, N540);
  nand NAND2_196 (N573, N488, N541);
  nand NAND2_197 (N577, N488, N542);
  nand NAND2_198 (N581, N488, N543);
  nand NAND2_204 (N590, N553, N159);
  nand NAND2_207 (N597, N557, N165);
  nand NAND2_210 (N606, N561, N171);
  nand NAND2_213 (N616, N565, N177);
  nand NAND2_216 (N625, N569, N183);
  nand NAND2_219 (N632, N573, N189);
  nand NAND2_222 (N641, N577, N195);
  nand NAND2_225 (N651, N581, N201);
  nand NAND2_254 (N732, N654, N261);
  nand NAND2_283 (N761, N644, N722);
  nand NAND2_284 (N762, N635, N713);
  nand NAND2_286 (N764, N609, N687);
  nand NAND2_287 (N765, N600, N678);
  nand NAND2_299 (N782, N651, N732);
  nand NAND2_310 (N795, N628, N773);
  nand NAND2_311 (N796, N795, N625);
  nand NAND2_322 (N812, N619, N796);
  nand NAND2_327 (N822, N616, N812);
  nand NAND2_344 (N841, N815, N593);
  nand NAND3_117 (N443, N447, N319, N17);
  nand NAND3_255 (N733, N644, N654, N261);
  nand NAND3_285 (N763, N635, N644, N722);
  nand NAND3_288 (N766, N600, N609, N687);
  nand NAND3_297 (N778, N641, N761, N733);
  nand NAND3_323 (N813, N609, N619, N796);
  nand NAND3_326 (N819, N606, N764, N813);
  nand NAND3_340 (N863, N826, N777, N704);
  nand NAND3_357 (N874, N845, N772, N696);
  nand NAND3_370 (N878, N859, N769, N669);
  nand NAND3_371 (N879, N860, N770, N677);
  nand NAND3_372 (N880, N861, N771, N686);
  nand NAND4_1 (N269, N1, N8, N13, N17);
  nand NAND4_2 (N270, N1, N26, N13, N17);
  nand NAND4_5 (N279, N1, N8, N51, N17);
  nand NAND4_6 (N280, N1, N8, N13, N55);
  nand NAND4_116 (N442, N375, N59, N156, N447);
  nand NAND4_256 (N734, N635, N644, N654, N261);
  nand NAND4_295 (N773, N632, N762, N763, N734);
  nand NAND4_321 (N850, N805, N787, N731, N529);
  nand NAND4_324 (N814, N600, N609, N619, N796);
  nand NAND4_325 (N815, N597, N765, N766, N814);
  nand NAND4_341 (N864, N827, N781, N712, N527);
  nand NAND4_342 (N865, N828, N785, N721, N528);
  nor NOR2_34 (N322, N17, N42);
  nor NOR2_74 (N375, N322, N323);
  nor NOR2_126 (N460, N406, N425);
  nor NOR2_127 (N463, N409, N426);
  nor NOR2_142 (N492, N413, N444);
  nor NOR2_143 (N495, N416, N445);
  nor NOR2_149 (N503, N475, N476);
  nor NOR2_151 (N505, N477, N476);
  nor NOR2_153 (N507, N479, N476);
  nor NOR2_155 (N509, N481, N476);
  nor NOR2_178 (N536, N309, N502);
  nor NOR2_179 (N537, N316, N504);
  nor NOR2_180 (N538, N317, N506);
  nor NOR2_181 (N539, N318, N508);
  nor NOR2_182 (N540, N510, N511);
  nor NOR2_183 (N541, N512, N513);
  nor NOR2_184 (N542, N514, N515);
  nor NOR2_185 (N543, N516, N517);
  nor NOR2_228 (N767, N552, N588);
  nor NOR2_229 (N768, N587, N589);
  nor NOR2_232 (N669, N596, N522);
  nor NOR2_235 (N677, N605, N523);
  nor NOR2_238 (N686, N615, N524);
  nor NOR2_241 (N696, N624, N525);
  nor NOR2_244 (N704, N631, N526);
  nor NOR2_247 (N712, N337, N640);
  nor NOR2_250 (N721, N339, N650);
  nor NOR2_253 (N731, N341, N659);
  nor NOR2_279 (N757, N727, N261);
  nor NOR2_291 (N769, N736, N737);
  nor NOR2_292 (N770, N739, N740);
  nor NOR2_293 (N771, N742, N743);
  nor NOR2_294 (N772, N745, N746);
  nor NOR2_296 (N777, N748, N749);
  nor NOR2_298 (N781, N751, N752);
  nor NOR2_300 (N785, N754, N755);
  nor NOR2_301 (N786, N757, N758);
  nor NOR2_302 (N787, N759, N760);
  nor NOR2_303 (N788, N700, N773);
  nor NOR2_305 (N790, N708, N778);
  nor NOR2_307 (N792, N717, N782);
  nor NOR2_312 (N802, N788, N789);
  nor NOR2_313 (N803, N790, N791);
  nor NOR2_314 (N804, N792, N793);
  nor NOR2_315 (N805, N340, N794);
  nor NOR2_316 (N806, N692, N796);
  nor NOR2_328 (N825, N806, N807);
  nor NOR2_329 (N826, N335, N808);
  nor NOR2_330 (N827, N336, N809);
  nor NOR2_331 (N828, N338, N810);
  nor NOR2_333 (N830, N665, N815);
  nor NOR2_335 (N832, N673, N819);
  nor NOR2_337 (N834, N682, N822);
  nor NOR2_345 (N842, N830, N831);
  nor NOR2_346 (N843, N832, N833);
  nor NOR2_347 (N844, N834, N835);
  nor NOR2_348 (N845, N334, N836);
  nor NOR2_362 (N859, N417, N851);
  nor NOR2_363 (N860, N332, N852);
  nor NOR2_364 (N861, N333, N853);
  not NOT1_54 (N418, N269);
  not NOT1_55 (N343, N390);
  not NOT1_59 (N347, N279);
  not NOT1_63 (N420, N293);
  not NOT1_64 (N352, N294);
  not NOT1_65 (N421, N295);
  not NOT1_66 (N422, N296);
  not NOT1_87 (N448, N349);
  not NOT1_88 (N449, N350);
  not NOT1_89 (N450, N355);
  not NOT1_90 (N404, N357);
  not NOT1_91 (N405, N360);
  not NOT1_93 (N407, N363);
  not NOT1_94 (N408, N366);
  not NOT1_97 (N411, N376);
  not NOT1_98 (N412, N379);
  not NOT1_100 (N414, N382);
  not NOT1_101 (N415, N385);
  not NOT1_188 (N550, N530);
  not NOT1_189 (N551, N533);
  not NOT1_199 (N585, N544);
  not NOT1_200 (N586, N547);
  not NOT1_230 (N662, N590);
  not NOT1_233 (N670, N597);
  not NOT1_236 (N678, N606);
  not NOT1_239 (N687, N616);
  not NOT1_242 (N697, N625);
  not NOT1_245 (N705, N632);
  not NOT1_248 (N713, N641);
  not NOT1_251 (N722, N651);
  not NOT1_361 (N866, N849);
  or OR2_19 (N298, N87, N88);
  or OR2_21 (N302, N91, N96);
  or OR2_23 (N304, N101, N106);
  or OR2_25 (N306, N111, N116);
  or OR2_27 (N308, N121, N126);
  or OR2_37 (N325, N159, N165);
  or OR2_39 (N327, N171, N177);
  or OR2_41 (N329, N183, N189);
  or OR2_43 (N331, N195, N201);
  or OR2_56 (N419, N270, N390);
  or OR2_61 (N349, N280, N285);
  or OR2_83 (N446, N270, N343);
  or OR2_145 (N499, N130, N460);
  or OR2_147 (N501, N463, N135);
  or OR2_165 (N519, N130, N492);
  or OR2_167 (N521, N495, N207);
  or OR2_205 (N593, N553, N159);
  or OR2_208 (N600, N557, N165);
  or OR2_211 (N609, N561, N171);
  or OR2_214 (N619, N565, N177);
  or OR2_217 (N628, N569, N183);
  or OR2_220 (N635, N573, N189);
  or OR2_223 (N644, N577, N195);
  or OR2_226 (N654, N581, N201);
  or g1 (N350, n_87, n_88, n_89, N280);
  not g2 (n_87, N59);
  not g3 (n_88, N68);
  not g4 (n_89, N74);
  and g5 (n_91, n_90, N59);
  not g6 (n_90, N280);
  and g7 (n_92, N42, N68);
  and g8 (N400, N72, N73, n_91, n_92);
  or g9 (N488, n_93, n_94, n_95, N268);
  not g10 (n_93, N447);
  not g11 (n_94, N287);
  not g12 (n_95, N55);
  and g13 (N476, n_96, N447, N17, N287);
  not g14 (n_96, N268);
endmodule